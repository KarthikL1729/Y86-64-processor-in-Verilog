module execute(clk)